module function_void;
function void welcome();
$display("==welcome==");
$display("==Hi==");
$display("==BY==");
endfunction
initial begin
welcome();
end
endmodule 
